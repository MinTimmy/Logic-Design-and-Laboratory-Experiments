library verilog;
use verilog.vl_types.all;
entity t_Moore_Model is
end t_Moore_Model;
