library verilog;
use verilog.vl_types.all;
entity Demo1_vlg_vec_tst is
end Demo1_vlg_vec_tst;
