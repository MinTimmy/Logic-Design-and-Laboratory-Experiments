library verilog;
use verilog.vl_types.all;
entity mux_4x1_beh_vlg_check_tst is
    port(
        m_out           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux_4x1_beh_vlg_check_tst;
