library verilog;
use verilog.vl_types.all;
entity JK_FF_vlg_check_tst is
    port(
        Q               : in     vl_logic;
        Q_b             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end JK_FF_vlg_check_tst;
