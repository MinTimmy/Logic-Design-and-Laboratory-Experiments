library verilog;
use verilog.vl_types.all;
entity Demo2_vlg_check_tst is
    port(
        m_out           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Demo2_vlg_check_tst;
