library verilog;
use verilog.vl_types.all;
entity test_Demo4 is
end test_Demo4;
