library verilog;
use verilog.vl_types.all;
entity Mealy_Zero_Detector_vlg_vec_tst is
end Mealy_Zero_Detector_vlg_vec_tst;
