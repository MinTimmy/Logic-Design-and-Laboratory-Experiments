library verilog;
use verilog.vl_types.all;
entity t_full_add is
end t_full_add;
