library verilog;
use verilog.vl_types.all;
entity t_Mealy_Zero_Detector is
end t_Mealy_Zero_Detector;
