library verilog;
use verilog.vl_types.all;
entity JK_Flip_flop_vlg_vec_tst is
end JK_Flip_flop_vlg_vec_tst;
