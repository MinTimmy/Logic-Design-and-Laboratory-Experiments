library verilog;
use verilog.vl_types.all;
entity D_Flip_flop_vlg_vec_tst is
end D_Flip_flop_vlg_vec_tst;
