library verilog;
use verilog.vl_types.all;
entity Demo2_vlg_vec_tst is
end Demo2_vlg_vec_tst;
